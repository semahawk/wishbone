`ifndef __PARAMETERS_SV__
`define __PARAMETERS_SV__

`define ADDR_WIDTH 8
`define DATA_WIDTH 8

`endif // __PARAMETERS_SV__
