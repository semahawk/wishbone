`ifndef __PARAMETERS_SV__
`define __PARAMETERS_SV__

`define ADDR_WIDTH 16
`define DATA_WIDTH 32

`endif // __PARAMETERS_SV__
